library verilog;
use verilog.vl_types.all;
entity tb_controller is
end tb_controller;
