library verilog;
use verilog.vl_types.all;
entity tb_Calculate_NTLM is
end tb_Calculate_NTLM;
