library verilog;
use verilog.vl_types.all;
entity tb_hashcracker is
end tb_hashcracker;
