// Code your testbench here
// or browse Examples
`timescale 1ns / 10ps

module tb_Calculate_NTLM_reg();
  
  parameter CLK_PERIOD				= 10;
  reg [0:127] tb_instr;
  reg [0:3] tb_length;
  reg [0:127] tb_hash;
  reg [0:127] tb_outstr;
  reg tb_clk;
  reg tb_n_rst;
  
  always
	begin : CLK_GEN
		tb_clk = 1'b0;
		#(CLK_PERIOD / 2);
		tb_clk = 1'b1;
		#(CLK_PERIOD / 2);
	end

	Calculate_NTLM_reg DUT
	(
   	.instr(tb_instr),
		.length(tb_length),
		.hash(tb_hash),
    .clk(tb_clk),
    .n_rst(tb_n_rst),
    .outstr(tb_outstr)
	);
	
	
	initial
	begin 
		 //tb_instr = 128'b01110000011000010111001101110011011101110110111100000000000000000000000000000000000000000000000000000000000000000000000000000000;
		 //tb_length = 6;
		 //tb_instr = 128'b01110000011000010111001101110011011101110110111101110010000000000000000000000000000000000000000000000000000000000000000000000000;
		 //tb_length = 7;
		 //tb_instr = 128'b01110000011000010111001101110011011101110110111101110010011001000000000000000000000000000000000000000000000000000000000000000000;
		 //tb_length = 8;
		 tb_instr[0:15] = 16'b0110001001100001;
		 tb_instr[16:127] = 0;
		 tb_length = 2;
		 tb_n_rst = 0;
    	#CLK_PERIOD
    	#1
    	tb_n_rst = 1;
    	//#CLK_PERIOD
    	//tb_instr = 128'b01100001011000010110000101100001011000010110000100000000000000000000000000000000000000000000000000000000000000000000000000000000;
		 //tb_length = 6;
    	//tb_instr = 128'b01110000011000010111001101110011011101110110111101110010000000000000000000000000000000000000000000000000000000000000000000000000;
		 //tb_length = 7;
		 //#CLK_PERIOD
		 //tb_instr = 128'b01100010011000010110001001100001011000100110000100000000000000000000000000000000000000000000000000000000000000000000000000000000;
		 //tb_length = 6;
    	//tb_instr = 128'b01110000011000010111001101110011011101110110111101110010011001000000000000000000000000000000000000000000000000000000000000000000;
		 //tb_length = 8;
 	
    end
endmodule