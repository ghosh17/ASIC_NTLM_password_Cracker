`timescale 1ns / 10ps
module Calculate_NTLM
(
    input wire [0:127] instr,
  	input wire [0:3] length,
    output reg [0:127] hash,
    output reg [0:511] buff,
  	//output reg [0:511] buff
  output reg [0:31] a4,
  output reg [0:31] b4,
  output reg [0:31] c4,
  output reg [0:31] d4
);
  reg [0:127] temphash;
	//reg [0:511] buff;
  parameter ai = 32'h67452301;
  parameter bi = 32'hefcdab89;
  parameter ci = 32'h98badcfe;
  parameter di = 32'h10325476;
  parameter root2 = 32'h5a827999;
  parameter root3 = 32'h6ed9eba1;
  reg [0:31] a1;
  reg [0:31] a2;
  reg [0:31] a3;
  //reg [0:31] a4;
  reg [0:31] a5;
  reg [0:31] a6;
  reg [0:31] a7;
  reg [0:31] a8;
  reg [0:31] a9;
  reg [0:31] a10;
  reg [0:31] a11;
  reg [0:31] a12;
  reg [0:31] a13;
  reg [0:31] a14;
  reg [0:31] a15;
  reg [0:31] a16;
  reg [0:31] a17;
  reg [0:31] a18;
  reg [0:31] a19;
  reg [0:31] a20;
  reg [0:31] a21;
  reg [0:31] a22;
  reg [0:31] a23;
  reg [0:31] a24;
  reg [0:31] b1;
  reg [0:31] b2;
  reg [0:31] b3;
  //reg [0:31] b4;
  reg [0:31] b5;
  reg [0:31] b6;
  reg [0:31] b7;
  reg [0:31] b8;
  reg [0:31] b9;
  reg [0:31] b10;
  reg [0:31] b11;
  reg [0:31] b12;
  reg [0:31] b13;
  reg [0:31] b14;
  reg [0:31] b15;
  reg [0:31] b16;
  reg [0:31] b17;
  reg [0:31] b18;
  reg [0:31] b19;
  reg [0:31] b20;
  reg [0:31] b21;
  reg [0:31] b22;
  reg [0:31] b23;
  reg [0:31] b24;
  reg [0:31] c1;
  reg [0:31] c2;
  reg [0:31] c3;
  //reg [0:31] c4;
  reg [0:31] c5;
  reg [0:31] c6;
  reg [0:31] c7;
  reg [0:31] c8;
  reg [0:31] c9;
  reg [0:31] c10;
  reg [0:31] c11;
  reg [0:31] c12;
  reg [0:31] c13;
  reg [0:31] c14;
  reg [0:31] c15;
  reg [0:31] c16;
  reg [0:31] c17;
  reg [0:31] c18;
  reg [0:31] c19;
  reg [0:31] c20;
  reg [0:31] c21;
  reg [0:31] c22;
  reg [0:31] c23;
  reg [0:31] c24;
  reg [0:31] d1;
  reg [0:31] d2;
  reg [0:31] d3;
  //reg [0:31] d4;
  reg [0:31] d5;
  reg [0:31] d6;
  reg [0:31] d7;
  reg [0:31] d8;
  reg [0:31] d9;
  reg [0:31] d10;
  reg [0:31] d11;
  reg [0:31] d12;
  reg [0:31] d13;
  reg [0:31] d14;
  reg [0:31] d15;
  reg [0:31] d16;
  reg [0:31] d17;
  reg [0:31] d18;
  reg [0:31] d19;
  reg [0:31] d20;
  reg [0:31] d21;
  reg [0:31] d22;
  reg [0:31] d23;
  reg [0:31] d24;
    always_comb 
        begin
          if(length >1)buff[32*0:32*0+31] = instr[2 * 8*0:2 * 8*0 +7] | (instr[8*(2 * 0 + 1):8*(2 * 0 + 1) + 7] << 16);//i=0
          if(length >3)buff[32*1:32*1+31] = instr[2 * 8*1:2 * 8*1 +7] | (instr[8*(2 * 1 + 1):8*(2 * 1 + 1) + 7] << 16);//i=1
          if(length >5)buff[32*2:32*2+31] = instr[2 * 8*2:2 * 8*2 +7] | (instr[8*(2 * 2 + 1):8*(2 * 2 + 1) + 7] << 16);//i=2
          if(length >7)buff[32*3:32*3+31] = instr[2 * 8*3:2 * 8*3 +7] | (instr[8*(2 * 3 + 1):8*(2 * 3 + 1) + 7] << 16);//i=3
          if(length >9)buff[32*4:32*4+31] = instr[2 * 8*4:2 * 8*4 +7] | (instr[8*(2 * 4 + 1):8*(2 * 4 + 1) + 7] << 16);//i=4
          if(length >11)buff[32*5:32*5+31] = instr[2 * 8*5:2 * 8*5 +7] | (instr[8*(2 * 5 + 1):8*(2 * 5 + 1) + 7] << 16);//i=5
          if(length >13)buff[32*6:32*6+31] = instr[2 * 8*6:2 * 8*6 +7] | (instr[8*(2 * 6 + 1):8*(2 * 6 + 1) + 7] << 16);//i=6
          if(length >15)buff[32*7:32*7+31] = instr[2 * 8*7:2 * 8*7 +7] | (instr[8*(2 * 7 + 1):8*(2 * 7 + 1) + 7] << 16);//i=7
          
          //padding
          if(length == 0) begin
            buff[32*(0/2):32*(0/2) + 31] = 8'h80;
            buff[32*(0/2) + 32:14*32 + 31] = length << 4;
          end
          else if(length == 1) begin
            buff[32*(1/2):32*(1/2) + 31] = instr[8*(1 - 1):8*(1 - 1) + 7] | 24'h800000;
            buff[32*(1/2) + 32:14*32 + 31] = length << 4;
            buff[15*32:15*32 + 31] = 0;
          end
          else if(length == 2)begin
            buff[32*(2/2):32*(2/2) + 31] = 8'h80;
            buff[32*(2/2) + 32:14*32 + 31] = length << 4;
            buff[15*32:15*32 + 31] = 0;
          end
          else if(length == 3) begin
            buff[32*(3/2):32*(3/2) + 31] = instr[8*(3 - 1):8*(3 - 1) + 7] | 24'h800000;
            buff[32*(3/2) + 32:14*32 + 31] = length << 4;
            buff[15*32:15*32 + 31] = 0;
          end
          else if(length == 4)begin
            buff[32*(4/2):32*(4/2) + 31] = 8'h80;
            buff[32*(4/2) + 32:14*32 + 31] = length << 4;
            buff[15*32:15*32 + 31] = 0;
          end
          else if(length == 5)begin
            buff[32*(5/2):32*(5/2) + 31] = instr[8*(5 - 1):8*(5 - 1) + 7] | 24'h800000;
            buff[32*(5/2) + 32:14*32 + 31] = length << 4;
            buff[15*32:15*32 + 31] = 0;
          end
          else if(length == 6)begin
            buff[32*(6/2):32*(6/2) + 31] = 8'h80;
            buff[32*(6/2) + 32:14*32 + 31] = length << 4;
            buff[15*32:15*32 + 31] = 0;
          end
          else if(length == 7)begin
            buff[32*(7/2):32*(7/2) + 31] = instr[8*(7 - 1):8*(7 - 1) + 7] | 24'h800000;
            buff[32*(7/2) + 32:14*32 + 31] = length << 4;
            buff[15*32:15*32 + 31] = 0;
          end
          else if(length == 8)begin
            buff[32*(8/2):32*(8/2) + 31] = 8'h80;
            buff[32*(8/2) + 32:14*32 + 31] = length << 4;
            buff[15*32:15*32 + 31] = 0;
          end
          else if(length == 9)begin
            buff[32*(9/2):32*(9/2) + 31] = instr[8*(9 - 1):8*(9 - 1) + 7] | 24'h800000;
            buff[32*(9/2) + 32:14*32 + 31] = length << 4;
            buff[15*32:15*32 + 31] = 0;
          end
          else if(length == 10)begin
            buff[32*(10/2):32*(10/2) + 31] = 8'h80;
            buff[32*(10/2) + 32:14*32 + 31] = length << 4;
            buff[15*32:15*32 + 31] = 0;
          end
          else if(length == 11)begin
            buff[32*(11/2):32*(11/2) + 31] = instr[8*(11 - 1):8*(11 - 1) + 7] | 24'h800000;
            buff[32*(11/2) + 32:14*32 + 31] = length << 4;
            buff[15*32:15*32 + 31] = 0;
          end
          else if(length == 12)begin
            buff[32*(12/2):32*(12/2) + 31] = 8'h80;
            buff[32*(12/2) + 32:14*32 + 31] = length << 4;
            buff[15*32:15*32 + 31] = 0;
          end
          else if(length == 13)begin
            buff[32*(13/2):32*(13/2) + 31] = instr[8*(13 - 1):8*(13 - 1) + 7] | 24'h800000;
            buff[32*(13/2) + 32:14*32 + 31] = length << 4;
            buff[15*32:15*32 + 31] = 0;
          end
          else if(length == 14)begin
            buff[32*(14/2):32*(14/2) + 31] = 8'h80;
            buff[32*(14/2) + 32:14*32 + 31] = length << 4;
            buff[15*32:15*32 + 31] = 0;
          end
          else if(length == 15)begin
            buff[32*(15/2):32*(15/2) + 31] = instr[8*(15 - 1):8*(15 - 1) + 7] | 24'h800000;
            buff[32*(15/2) + 32:14*32 + 31] = length << 4;
            buff[15*32:15*32 + 31] = 0;
          end
          else begin//Length 16, realistically it should not get higher than this (avoiding a latch here)
            buff[32*(16/2):32*(16/2) + 31] = 8'h80;
            buff[32*(16/2) + 32:14*32 + 31] = length << 4;
            buff[15*32:15*32 + 31] = 0;
          end
		  
          //put the length
          //buff[14*32:14*32 + 31] = length << 4;
          /* Round 1 */
          a1 = ai + ((di ^ (bi & (ci ^ di)))  +  buff[32*0 : 32*0 + 31]);
          a2 = (a1 << 3 ) | (a1 >> 29);
          d1 = di + ((ci ^ (a2 & (bi ^ ci)))  +  buff[32*1 : 32*1 + 31]);
          d2 = (d1 << 7 ) | (d1 >> 25);
          c1 = ci + ((bi ^ (d2 & (a2 ^ bi)))  +  buff[2*32 : 2*32 + 31]);
          c2 = (c1 << 11) | (c1 >> 21);
          b1 = bi + ((a2 ^ (c2 & (d2 ^ a2)))  +  buff[3*32 : 3*32 + 31]);
          b2 = (b1 << 19) | (b1 >> 13);
          
          a3 = a2 + ((d2 ^ (b2 & (c2 ^ d2)))  +  buff[32*4 : 32*4 + 31])  ;
          a4 = (a3 << 3 ) | (a3 >> 29);
          d3 = d2 + ((c2 ^ (a4 & (b2 ^ c2)))  +  buff[32*5 : 32*5 + 31])  ;
          d4 = (d3 << 7 ) | (d3 >> 25);
          c3 = c2 + ((b2 ^ (d4 & (a4 ^ b2)))  +  buff[32*6 : 32*6 + 31])  ;
          c4 = (c3 << 11) | (c3 >> 21);
          b3 = b2 + ((a4 ^ (c4 & (d4 ^ a4)))  +  buff[32*7 : 32*7 + 31])  ;
          b4 = (b3 << 19) | (b3 >> 13);
 
          a5 = a4 + ((d4 ^ (b4 & (c4 ^ d4)))  +  buff[32*8 : 32*8 + 31])  ;
          a6 = (a5 << 3 ) | (a5 >> 29);
          d5 = d4 + ((c4 ^ (a6 & (b4 ^ c4)))  +  buff[32*9 : 32*9 + 31]) ;
          d6 = (d5 << 7 ) | (d5 >> 25);
          c5 = c4 + ((b4 ^ (d6 & (a6 ^ b4)))  +  buff[32*10 : 32*10 + 31]) ;
          c6 = (c5 << 11) | (c5 >> 21);
          b5 = b4 + ((a6 ^ (c6 & (d6 ^ a6)))  +  buff[32*11 : 32*11 + 31]) ;
          b6 = (b5 << 19) | (b5 >> 13);
 
          a7 = a6 + (d6 ^ (b6 & (c6 ^ d6)))  +  buff[32*12 : 32*12 + 31] ;
          a8 = (a7 << 3 ) | (a7 >> 29);
          d7 = d6 + (c6 ^ (a8 & (b6 ^ c6)))  +  buff[32*13 : 32*13 + 31] ;
          d8 = (d7 << 7 ) | (d7 >> 25);
          c7 = c6 + (b6 ^ (d8 & (a8 ^ b6)))  +  buff[32*14 : 32*14 + 31] ;
          c8 = (c7 << 11) | (c7 >> 21);
          b7 = b6 + (a8 ^ (c8 & (d8 ^ a8)))  +  buff[32*15 : 32*15 + 31] ;
          b8 = (b7 << 19) | (b7 >> 13);
 
	/* Round 2 */
          a9 = a8 + ((b8 & (c8 | d8)) | (c8 & d8)) + buff[32*0 : 32*0 + 31] +root2; 
          a10 = (a9<<3 ) | (a9>>29);
          d9 = d8 + ((a10 & (b8 | c8)) | (b8 & c8)) + buff[32*4 : 32*4 + 31] +root2; 
          d10 = (d9<<5 ) | (d9>>27);
          c9 = c8 + ((d10 & (a10 | b8)) | (a10 & b8)) + buff[32*8 : 32*8 + 31] +root2; 
          c10 = (c9<<9 ) | (c9>>23);
          b9 = b8 + ((c10 & (d10 | a10)) | (d10 & a10)) + buff[32*12 : 32*12 + 31]+root2; 
          b10 = (b9<<13) | (b9>>19);
 
          a11 = a10 + ((b10 & (c10 | d10)) | (c10 & d10)) + buff[32*1 : 32*1 + 31] +root2; 
          a12 = (a11<<3 ) | (a11>>29);
          d11 = d10 + ((a12 & (b10 | c10)) | (b10 & c10)) + buff[32*5 : 32*5 + 31] +root2; 
          d12 = (d11<<5 ) | (d11>>27);
          c11 = c10 + ((d12 & (a12 | b10)) | (a12 & b10)) + buff[32*9 : 32*9 + 31] +root2; 
          c12 = (c11<<9 ) | (c11>>23);
          b11 = b10 + ((c12 & (d12 | a12)) | (d12 & a12)) + buff[32*13 : 32*13 + 31]+root2; 
          b12 = (b11<<13) | (b11>>19);
 
          a13 = a12 + ((b12 & (c12 | d12)) | (c12 & d12)) + buff[32*2 : 32*2 + 31] +root2; 
          a14 = (a13<<3 ) | (a13>>29);
          d13 = d12 + ((a14 & (b12 | c12)) | (b12 & c12)) + buff[32*6 : 32*6 + 31] +root2; 
          d14 = (d13<<5 ) | (d13>>27);
          c13 = c12 +((d14 & (a14 | b12)) | (a14 & b12)) + buff[32*10 : 32*10 + 31]+root2; 
          c14 = (c13<<9 ) | (c13>>23);
          b13 = b12 + ((c14 & (d14 | a14)) | (d14 & a14)) + buff[32*14 : 32*14 + 31]+root2; 
          b14 = (b13<<13) | (b13>>19);
 
          a15 = a14 + ((b14 & (c14 | d14)) | (c14 & d14)) + buff[32*3 : 32*3 + 31] +root2; 
          a16 = (a15<<3 ) | (a15>>29);
          d15 = d14 + ((a16 & (b14 | c14)) | (b14 & c14)) + buff[32*7 : 32*7 + 31] +root2; 
          d16 = (d15<<5 ) | (d15>>27);
          c15 = c14 + ((d16 & (a16 | b14)) | (a16 & b14)) + buff[32*11 : 32*11 + 31]+root2; 
          c16 = (c15<<9 ) | (c15>>23);
          b15 = b14 + ((c16 & (d16 | a16)) | (d16 & a16)) + buff[32*15 : 32*15 + 31]+root2; 
          b16 = (b15<<13) | (b15>>19);
 
	/* Round 3 */
          a17 = a16 + (d16 ^ c16 ^ b16) + buff[32*0 : 32*0 + 31]  +  root3; 
          a18 = (a17 << 3 ) | (a17 >> 29);
          d17 = d16 + (c16 ^ b16 ^ a18) + buff[32*8 : 32*8 + 31]  +  root3; 
          d18 = (d17 << 9 ) | (d17 >> 23);
          c17 = c16 + (b16 ^ a18 ^ d18) + buff[32*4 : 32*4 + 31]  +  root3; 
          c18 = (c17 << 11) | (c17 >> 21);
          b17 = b16 + (a18 ^ d18 ^ c18) + buff[32*12 : 32*12 + 31] +  root3; 
          b18 = (b17 << 15) | (b17 >> 17);
 
          a19 = a18 + (d18 ^ c18 ^ b18) + buff[32*2 : 32*2 + 31]  +  root3; 
          a20 = (a19 << 3 ) | (a19 >> 29);
          d19 = d18 + (c18 ^ b18 ^ a20) + buff[32*10 : 32*10 + 31] +  root3; 
          d20 = (d19 << 9 ) | (d19 >> 23);
          c19 = c18 + (b18 ^ a20 ^ d20) + buff[32*6 : 32*6 + 31]  +  root3; 
          c20 = (c19 << 11) | (c19 >> 21);
          b19 = b18 + (a20 ^ d20 ^ c20) + buff[32*14 : 32*14 + 31] +  root3; 
          b20 = (b19 << 15) | (b19 >> 17);
 
          a21 = a20 + (d20 ^ c20 ^ b20) + buff[32*1 : 32*1 + 31]  +  root3; 
          a22 = (a21 << 3 ) | (a21 >> 29);
          d21 = d20 + (c20 ^ b20 ^ a22) + buff[32*9 : 32*9 + 31]  +  root3; 
          d22 = (d21 << 9 ) | (d21 >> 23);
          c21 = c20 + (b20 ^ a22 ^ d22) + buff[32*5 : 32*5 + 31]  +  root3; 
          c22 = (c21 << 11) | (c21 >> 21);
          b21 = b20 + (a22 ^ d22 ^ c22) + buff[32*13 : 32*13 + 31] +  root3; 
          b22 = (b21 << 15) | (b21 >> 17);
 
          a23 = a22 + (d22 ^ c22 ^ b22) + buff[32*3 : 32*3 + 31]  +  root3; 
          a24 = (a23 << 3 ) | (a23 >> 29);
          d23 = d22 + (c22 ^ b22 ^ a24) + buff[32*11 : 32*11 + 31] +  root3; 
          d24 = (d23 << 9 ) | (d23 >> 23);
          c23 = c22 + (b22 ^ a24 ^ d24) + buff[32*7 : 32*7 + 31]  +  root3; 
          c24 = (c23 << 11) | (c23 >> 21);
          b23 = b22 + (a24 ^ d24 ^ c24) + buff[32*15 : 32*15 + 31] +  root3; 
          b24 = (b23 << 15) | (b23 >> 17);
 
          temphash[0:31] = a24 + ai;
          temphash[32:63] = b24 + bi;
          temphash[64:95] = c24 + ci;
          temphash[96:127] = d24 + di;
          
          hash[0*8:1*8 - 1] = temphash[3*8:4*8 - 1];
          hash[1*8:2*8 - 1] = temphash[2*8:3*8 - 1];
          hash[2*8:3*8 - 1] = temphash[1*8:2*8 - 1];
          hash[3*8:4*8 - 1] = temphash[0*8:1*8 - 1];
          
          hash[4*8:5*8 - 1] = temphash[7*8:8*8 - 1];
          hash[5*8:6*8 - 1] = temphash[6*8:7*8 - 1];
          hash[6*8:7*8 - 1] = temphash[5*8:6*8 - 1];
          hash[7*8:8*8 - 1] = temphash[4*8:5*8 - 1];
          
          hash[8*8:9*8 - 1] = temphash[11*8:12*8 - 1];
          hash[9*8:10*8 - 1] = temphash[10*8:11*8 - 1];
          hash[10*8:11*8 - 1] = temphash[9*8:10*8 - 1];
          hash[11*8:12*8 - 1] = temphash[8*8:9*8 - 1];
          
          hash[12*8:13*8 - 1] = temphash[15*8:16*8 - 1];
          hash[13*8:14*8 - 1] = temphash[14*8:15*8 - 1];
          hash[14*8:15*8 - 1] = temphash[13*8:14*8 - 1];
          hash[15*8:16*8 - 1] = temphash[12*8:13*8 - 1];
        end
endmodule
